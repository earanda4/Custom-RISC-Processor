// Code your testbench here
// or browse Examples
//`include "new_fix2flt_tb.sv"
`include "flt2fix_tb.sv"